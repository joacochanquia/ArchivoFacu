library verilog;
use verilog.vl_types.all;
entity DiagCont60 is
    port(
        C               : out    vl_logic;
        CLK             : in     vl_logic
    );
end DiagCont60;

library verilog;
use verilog.vl_types.all;
entity Prueba1 is
    port(
        D               : out    vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : out    vl_logic
    );
end Prueba1;

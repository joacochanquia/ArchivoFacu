library verilog;
use verilog.vl_types.all;
entity LatchNAND_vlg_vec_tst is
end LatchNAND_vlg_vec_tst;

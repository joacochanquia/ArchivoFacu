library verilog;
use verilog.vl_types.all;
entity GenPar_vlg_vec_tst is
end GenPar_vlg_vec_tst;

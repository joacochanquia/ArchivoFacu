library verilog;
use verilog.vl_types.all;
entity GenQ0_vlg_check_tst is
    port(
        Q0m             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end GenQ0_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity GenQ2_vlg_check_tst is
    port(
        Q2m             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end GenQ2_vlg_check_tst;

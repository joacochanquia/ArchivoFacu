library verilog;
use verilog.vl_types.all;
entity Flags_vlg_vec_tst is
end Flags_vlg_vec_tst;

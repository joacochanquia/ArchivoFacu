library verilog;
use verilog.vl_types.all;
entity MaquinaMoore_vlg_vec_tst is
end MaquinaMoore_vlg_vec_tst;

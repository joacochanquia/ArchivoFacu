library verilog;
use verilog.vl_types.all;
entity GenQ1_vlg_vec_tst is
end GenQ1_vlg_vec_tst;

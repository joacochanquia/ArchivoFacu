library verilog;
use verilog.vl_types.all;
entity Resta_vlg_vec_tst is
end Resta_vlg_vec_tst;

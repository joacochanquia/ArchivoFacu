library verilog;
use verilog.vl_types.all;
entity AND4b_vlg_vec_tst is
end AND4b_vlg_vec_tst;

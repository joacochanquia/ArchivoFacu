library verilog;
use verilog.vl_types.all;
entity DiagCont5_vlg_vec_tst is
end DiagCont5_vlg_vec_tst;

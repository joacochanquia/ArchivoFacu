library verilog;
use verilog.vl_types.all;
entity OR4b_vlg_vec_tst is
end OR4b_vlg_vec_tst;

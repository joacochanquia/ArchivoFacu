library verilog;
use verilog.vl_types.all;
entity DiagCont3_vlg_vec_tst is
end DiagCont3_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity DiagCont60_vlg_vec_tst is
end DiagCont60_vlg_vec_tst;

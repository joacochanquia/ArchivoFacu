library verilog;
use verilog.vl_types.all;
entity GeneradorEstado_vlg_vec_tst is
end GeneradorEstado_vlg_vec_tst;

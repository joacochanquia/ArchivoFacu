library verilog;
use verilog.vl_types.all;
entity DetMagRel1bit_vlg_vec_tst is
end DetMagRel1bit_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity GenQ1_vlg_check_tst is
    port(
        Q1m             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end GenQ1_vlg_check_tst;

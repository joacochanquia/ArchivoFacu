library verilog;
use verilog.vl_types.all;
entity INC_vlg_vec_tst is
end INC_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity CA2_vlg_vec_tst is
end CA2_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity DiagCont3_vlg_check_tst is
    port(
        C               : in     vl_logic;
        Q0              : in     vl_logic;
        Q1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end DiagCont3_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity Flags_vlg_check_tst is
    port(
        N               : in     vl_logic;
        Z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Flags_vlg_check_tst;

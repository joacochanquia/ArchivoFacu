library verilog;
use verilog.vl_types.all;
entity MaquinaMoore2_vlg_vec_tst is
end MaquinaMoore2_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity GeneradorSalidas_vlg_vec_tst is
end GeneradorSalidas_vlg_vec_tst;

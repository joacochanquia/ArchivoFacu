library verilog;
use verilog.vl_types.all;
entity DiagCont3_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end DiagCont3_vlg_sample_tst;

library verilog;
use verilog.vl_types.all;
entity LatchNOR_vlg_vec_tst is
end LatchNOR_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Sumador2bits_vlg_vec_tst is
end Sumador2bits_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity GenQ3_vlg_check_tst is
    port(
        Q3m             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end GenQ3_vlg_check_tst;

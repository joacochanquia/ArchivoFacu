library verilog;
use verilog.vl_types.all;
entity XOR4b_vlg_vec_tst is
end XOR4b_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity DiagCont2_vlg_vec_tst is
end DiagCont2_vlg_vec_tst;

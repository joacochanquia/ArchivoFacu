library verilog;
use verilog.vl_types.all;
entity DetPar_vlg_vec_tst is
end DetPar_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity DecOp_vlg_vec_tst is
end DecOp_vlg_vec_tst;

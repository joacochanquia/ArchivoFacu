library verilog;
use verilog.vl_types.all;
entity GenQ0_vlg_vec_tst is
end GenQ0_vlg_vec_tst;

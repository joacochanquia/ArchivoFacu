library verilog;
use verilog.vl_types.all;
entity Suma_vlg_vec_tst is
end Suma_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity GenQ3_vlg_vec_tst is
end GenQ3_vlg_vec_tst;

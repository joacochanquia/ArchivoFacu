library verilog;
use verilog.vl_types.all;
entity Prueba1_vlg_vec_tst is
end Prueba1_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity BufferRetrasador_vlg_vec_tst is
end BufferRetrasador_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity SumaResta_vlg_vec_tst is
end SumaResta_vlg_vec_tst;

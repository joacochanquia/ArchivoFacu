library verilog;
use verilog.vl_types.all;
entity MaquinaMoore2_vlg_sample_tst is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        CLK             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end MaquinaMoore2_vlg_sample_tst;

library verilog;
use verilog.vl_types.all;
entity ABALU_vlg_vec_tst is
end ABALU_vlg_vec_tst;

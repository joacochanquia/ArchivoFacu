library verilog;
use verilog.vl_types.all;
entity DetMagRel3bit_vlg_check_tst is
    port(
        M               : in     vl_logic;
        N               : in     vl_logic;
        P               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end DetMagRel3bit_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity DiagCont2_vlg_check_tst is
    port(
        C               : in     vl_logic;
        Q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end DiagCont2_vlg_check_tst;

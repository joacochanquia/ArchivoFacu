library verilog;
use verilog.vl_types.all;
entity DetMagRel3bit_vlg_vec_tst is
end DetMagRel3bit_vlg_vec_tst;

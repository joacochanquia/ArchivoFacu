library verilog;
use verilog.vl_types.all;
entity GenQ2_vlg_vec_tst is
end GenQ2_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity BufferRetrasador_vlg_sample_tst is
    port(
        E               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end BufferRetrasador_vlg_sample_tst;

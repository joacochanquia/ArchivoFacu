library verilog;
use verilog.vl_types.all;
entity RegistroA_vlg_vec_tst is
end RegistroA_vlg_vec_tst;
